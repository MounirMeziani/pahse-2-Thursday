
library IEEE;
use ieee.std_logic_1164.all;

ENTITY con_ff_logic_tb IS
END;

ARCHITECTURE con_ff_logic_tb_arch of con_ff_logic_tb IS

signal busmuxin_TB :  STD_LOGIC_VECTOR(31 downto 0);
signal IRin_TB		 :  STD_LOGIC_VECTOR(1 downto 0);
signal CONin_TB 	 :  STD_LOGIC;
signal O_TB			 :  STD_LOGIC;
signal CLK         :  STD_LOGIC;
COMPONENT con_ff_logic
		PORT  (
			busmuxin	: IN STD_LOGIC_VECTOR(31 downto 0);
			IRin		: IN STD_LOGIC_VECTOR(1 downto 0);
			CONin 	: IN STD_LOGIC;
			O			: OUT STD_LOGIC
			);
END COMPONENT con_ff_logic;
	
BEGIN
	
	DUT1 : con_ff_logic
	
	PORT MAP (
		busmuxin => busmuxin_TB,
		IRin => IRin_TB,
		CONin => CONin_TB,
		O => O_TB
		
		);
		
	Clock_process: PROCESS
		BEGIN
			CLK <= '1', '0' after 10 ns;
			wait for 20 ns;
		END PROCESS CLK;
		
	process
	begin
	
		busmuxin <= b"11110000000000001111000000000000";
		
		
		IRin_TB <= b"00";
		IRin_TB <= b"01" after 40 ns;
		IRin_TB <= b"10" after 80 ns;
		IRin_TB <= b"11" after 120 ns;
		CONin_TB <= '1', '0' after 160 ns;
		
		wait;
	
	end process;
	
	end;